----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    02:05:37 02/18/2019 
-- Design Name: 
-- Module Name:    OR32BIT - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity OR32BIT is
    Port ( ORA : in  STD_LOGIC_VECTOR (31 downto 0);
           ORB : in  STD_LOGIC_VECTOR (31 downto 0);
           OROUT : out  STD_LOGIC_VECTOR (31 downto 0));
end OR32BIT;

architecture Behavioral of OR32BIT is

begin

OROUT <= ORA OR ORB AFTER 10 NS;

end Behavioral;

