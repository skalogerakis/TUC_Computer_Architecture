--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   22:32:11 02/20/2019
-- Design Name:   
-- Module Name:   C:/Xilinx/lab1_B/decoder5x32_TEST.vhd
-- Project Name:  lab1_B
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: decoder5x32
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY decoder5x32_TEST IS
END decoder5x32_TEST;
 
ARCHITECTURE behavior OF decoder5x32_TEST IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT decoder5x32
    PORT(
         decIN : IN  std_logic_vector(4 downto 0);
         decOUT : OUT  std_logic_vector(31 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal decIN : std_logic_vector(4 downto 0) := (others => '0');

 	--Outputs
   signal decOUT : std_logic_vector(31 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
   
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: decoder5x32 PORT MAP (
          decIN => decIN,
          decOUT => decOUT
        );

   -- Clock process definitions
  

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		
		
		
      decIN <="01100";
		wait for 100 ns;	
		
		decIN <="11111";
		wait for 100 ns;	
		
		decIN <="11000";
		wait for 100 ns;	
     
	   
	   
      -- insert stimulus here 

      wait;
   end process;

END;
