----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    19:56:49 03/14/2019 
-- Design Name: 
-- Module Name:    shiftBox - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity shiftBox is
			port (
			imm32_in: in std_logic_vector(31 downto 0);
			OpCode: in std_logic;
			imm32_out: out std_logic_vector(31 downto 0)
			);
end shiftBox;
			
architecture Behavioral of shiftBox is

begin

process(OpCode,imm32_in)
	
begin
	
	if (OpCode='1') then
	
	imm32_out <= imm32_in(29 downto 0) & "00";
	
	else 
	imm32_out <= imm32_in ;
	
	end if;

end process;

end Behavioral;

